module if_id.sv();

endmodule